`timescale 1ns / 1ps

module data_mem(
    input               clk, 
    input               mem_read_in,
    input               mem_write_in,
    input       [63:0]  alu_result_in,
    input       [63:0]  rs2_data_in,
    output reg  [63:0]  mem_read_data,
	output reg  [11:0]  addr_out
);
    wire [11:0] bram_addr = alu_result_in[11:0]; 
    reg [63:0] memory [0:4095];
    wire bram_en = mem_read_in | mem_write_in;
    wire bram_we = mem_write_in;
		initial begin: init_data_mem
        integer i;
        // 先將整塊記憶體清空為 0
        for(i = 0; i < 200; i = i + 1) begin
            memory[i] = 64'd0;
        end

        // ---------------------------------------------------------
        // 1. Vector Add 測試資料 (Int16)
        // 陣列 A 放 addr 0, 陣列 B 放 addr 1, 運算結果 C 預計存入 addr 2
        // ---------------------------------------------------------
        // A = {4, 3, 2, 1}
        memory[0] = 64'h0004_0003_0002_0001; 
        // B = {40, 30, 20, 10}
        memory[1] = 64'h0028_001E_0014_000A; 
        // [預期結果存於 addr 2] C = {44, 33, 22, 11} -> 64'h002C_0021_0016_000B

        // ---------------------------------------------------------
        // 2. Vector Sub 測試資料 (Int16)
        // 陣列 A 放 addr 10, 陣列 B 放 addr 11, 運算結果 C 預計存入 addr 12
        // ---------------------------------------------------------
        // A = {40, 30, 20, 10}
        memory[10] = 64'h0028_001E_0014_000A;
        // B = {4, 3, 2, 1}
        memory[11] = 64'h0004_0003_0002_0001;
        // [預期結果存於 addr 12] C = {36, 27, 18, 9} -> 64'h0024_001B_0012_0009

        // ---------------------------------------------------------
        // 3. BFloat16 向量乘法測試資料 (BF16)
        // 陣列 A 放 addr 20, 陣列 B 放 addr 21, 運算結果 C 預計存入 addr 22
        // BFloat16 格式參考: 1.0=3F80, 2.0=4000, 3.0=4040, -2.0=C000
        // ---------------------------------------------------------
        // A = {1.0, -2.0, 3.0, 2.0} 
        memory[20] = 64'h3F80_C000_4040_4000;
        // B = {2.0,  2.0, 2.0, 3.0}
        memory[21] = 64'h4000_4000_4000_4040;
        // [預期結果存於 addr 22] C = {2.0, -4.0, 6.0, 6.0} -> 64'h4000_C080_40C0_40C0

        // ---------------------------------------------------------
        // 4. BFloat16 融合乘加 (FMA) 測試資料 (BF16)
        // A 放 addr 30, B 放 addr 31, C 放 addr 32, 結果 D 存入 addr 33
        // ---------------------------------------------------------
        // A = {2.0, 2.0, 2.0, 2.0}
        memory[30] = 64'h4000_4000_4000_4000;
        // B = {3.0, 3.0, 3.0, 3.0}
        memory[31] = 64'h4040_4040_4040_4040;
        // C = {1.0, 1.0, 1.0, 1.0}
        memory[32] = 64'h3F80_3F80_3F80_3F80;
        // [預期結果存於 addr 33] D = A*B+C = {7.0, 7.0, 7.0, 7.0} -> 64'h40E0_40E0_40E0_40E0

        // ---------------------------------------------------------
        // 5. ReLU 激勵函數測試資料 (Int16)
        // 輸入 In 放 addr 40, 運算結果 Out 預計存入 addr 41
        // (複數以 2's complement 表示: -3=FFFD, -5=FFFB)
        // ---------------------------------------------------------
        // In = {8, -3, 10, -5}
        memory[40] = 64'h0008_FFFD_000A_FFFB;
        // [預期結果存於 addr 41] Out = max(0, In) = {8, 0, 10, 0} -> 64'h0008_0000_000A_0000
        
        // --- 設定記憶體推進常數 ---
        // 把數字 1 放在記憶體最後面，方便你的機器碼讀進 r10 當作推進指標的步長 (ADDI的替代品)
        //memory[4095] = 64'h0000_0000_0000_0001; 
    end
    always @(posedge clk) begin
        if (bram_en) begin
            if (bram_we) begin
                memory[bram_addr] <= rs2_data_in;
            end
            mem_read_data <= memory[bram_addr];
        end
    end
	
	always@(posedge clk)begin
		if (bram_en) begin
            addr_out <= bram_addr;
        end
	end
endmodule